`define TIMER_ADDR_W 2  //address width
`define TIMER_WDATA_W 1 //write data width
`define TIMER_RDATA_W 32//read data witdh
`ifndef DATA_W
 `define DATA_W 32      //cpu data width
`endif
